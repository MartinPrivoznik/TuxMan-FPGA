--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 


library IEEE;
use IEEE.STD_LOGIC_1164.all;

package ROM_Textures is

type square_resolution is array (0 to 15, 0 to 15) of STD_LOGIC_VECTOR(7 downto 0); -- RRRGGGBB

constant wall_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011")),
(("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"),("00000011"))
);

constant tuxman_closed_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000")),
(("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant tuxman_open_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant point_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111111"),("11111111"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111111"),("11111111"),("11111111"),("11111111"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111111"),("11111111"),("11111111"),("11111111"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111111"),("11111111"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant redghost_open_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"))
);
 
constant redghost_closed_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000")),
(("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("11100000"),("11100000"),("11100000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11100000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant blueghost_open_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"))
);
 
constant blueghost_closed_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011")),
(("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00011011"),("00011011"),("00011011"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00011011"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant greenghost_open_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101")),
(("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"))
);
 
constant greenghost_closed_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101")),
(("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101")),
(("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("10011101"),("10011101"),("10011101"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("10011101"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant yellowghost_open_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100")),
(("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"))
);
 
constant yellowghost_closed_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100")),
(("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100")),
(("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("11111100"),("11111100"),("11111100"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("11111100"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000")),
(("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"),("00000000"))
);

constant textblock_texture : Square_Resolution := 
(--  0             1            2            3            4            5            6            7            8            9            10           11           12           13          14           15
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111")),
(("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"),("11111111"))
);

end ROM_Textures;
